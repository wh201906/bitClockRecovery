
module globalClock (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
